//-------------------------------------------------------------------------
//						mem_sequencer - www.verificationguide.com
//-------------------------------------------------------------------------

class mem_sequencer extends uvm_sequencer#(mem_sequence_item);

    `uvm_component_utils(mem_sequencer) 
  
    //---------------------------------------
    //constructor
    //---------------------------------------
    function new(string name, uvm_component parent);
      super.new(name,parent);
    endfunction
    
  endclass